/nethome/amojumdar6/New_DV_Onboarding_Abhik/src/verilog/calc_tb_pkg.sv