/nethome/amojumdar6/New_DV_Onboarding_Abhik/src/verilog/result_buffer.sv