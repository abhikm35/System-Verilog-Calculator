/nethome/amojumdar6/New_DV_Onboarding_Abhik/src/verilog/full_adder.sv